----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:38:03 04/07/2014 
-- Design Name: 
-- Module Name:    Decoder32 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Decoder32 is
    Port ( I : in  STD_LOGIC_VECTOR (4 downto 0);
           O : out STD_LOGIC_VECTOR (31 downto 0);
           E : in  STD_LOGIC);
end Decoder32;

architecture Behavioral of Decoder32 is

begin
	O <= "00000000000000000000000000000000" WHEN E= '0' ELSE
	"00000000000000000000000000000001" WHEN I= "00000" ELSE
	"00000000000000000000000000000010" WHEN I= "00001" ELSE
	"00000000000000000000000000000100" WHEN I= "00010" ELSE
	"00000000000000000000000000001000" WHEN I= "00011" ELSE
	"00000000000000000000000000010000" WHEN I= "00100" ELSE
	"00000000000000000000000000100000" WHEN I= "00101" ELSE
	"00000000000000000000000001000000" WHEN I= "00110" ELSE
	"00000000000000000000000010000000" WHEN I= "00111" ELSE
	"00000000000000000000000100000000" WHEN I= "01000" ELSE
	"00000000000000000000001000000000" WHEN I= "01001" ELSE
	"00000000000000000000010000000000" WHEN I= "01010" ELSE
	"00000000000000000000100000000000" WHEN I= "01011" ELSE
	"00000000000000000001000000000000" WHEN I= "01100" ELSE
	"00000000000000000010000000000000" WHEN I= "01101" ELSE
	"00000000000000000100000000000000" WHEN I= "01110" ELSE
	"00000000000000001000000000000000" WHEN I= "01111" ELSE
	"00000000000000010000000000000000" WHEN I= "10000" ELSE
	"00000000000000100000000000000000" WHEN I= "10001" ELSE
	"00000000000001000000000000000000" WHEN I= "10010" ELSE
	"00000000000010000000000000000000" WHEN I= "10011" ELSE
	"00000000000100000000000000000000" WHEN I= "10100" ELSE
	"00000000001000000000000000000000" WHEN I= "10101" ELSE
	"00000000010000000000000000000000" WHEN I= "10110" ELSE
	"00000000100000000000000000000000" WHEN I= "10111" ELSE
	"00000001000000000000000000000000" WHEN I= "11000" ELSE
	"00000010000000000000000000000000" WHEN I= "11001" ELSE
	"00000100000000000000000000000000" WHEN I= "11010" ELSE
	"00001000000000000000000000000000" WHEN I= "11011" ELSE
	"00010000000000000000000000000000" WHEN I= "11100" ELSE
	"00100000000000000000000000000000" WHEN I= "11101" ELSE
	"01000000000000000000000000000000" WHEN I= "11110" ELSE
	"10000000000000000000000000000000" WHEN I= "11111" ELSE
	"XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX" ;
end Behavioral;

